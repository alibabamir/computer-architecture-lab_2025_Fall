 
--
----------------------------------------------------------------------------------
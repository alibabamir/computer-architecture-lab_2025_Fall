library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity tb_ripple_counter_tff is
    -- Testbench has no ports
end tb_ripple_counter_tff;

architecture Behavioral of tb_ripple_counter_tff is
    -- Component declaration for the ripple counter
    component ripple_counter_tff
        Port (
            clk     : in  STD_LOGIC;
            reset_n : in  STD_LOGIC;
            q       : out STD_LOGIC_VECTOR(3 downto 0)
        );
    end component;

    -- Testbench signals
    signal clk     : STD_LOGIC := '0';
    signal reset_n : STD_LOGIC := '1';
    signal q       : STD_LOGIC_VECTOR(3 downto 0);

    -- Clock period constant
    constant clk_period : time := 1 ns;

begin
    -- Instantiate the ripple counter
    uut: ripple_counter_tff
        Port map (
            clk     => clk,
            reset_n => reset_n,
            q       => q
        );

    -- Clock generation process
    clk_process: process
    begin
        clk <= '0';
        wait for clk_period / 2;
        clk <= '1';
        wait for clk_period / 2;
    end process;

    -- Stimulus process
    stimulus_process: process
    begin
        -- Apply reset
        reset_n <= '0';    -- Assert reset
        wait for 20 ns;
        reset_n <= '1';    -- Deassert reset
        wait for 100 ns;   -- Observe counter behavior

        -- Apply another reset after some time
        wait for 50 ns;
        reset_n <= '0';
        wait for 20 ns;
        reset_n <= '1';
        wait for 100 ns;

        -- End of simulation
        wait;
    end process;
end Behavioral;